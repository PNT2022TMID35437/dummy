// Actel Corporation Proprietary and Confidential
//  Copyright 2008 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
//  Revision Information:
// Jun09    Revision 4.1
// Aug10    Revision 4.2
// SVN Revision Information:
// SVN $Revision: 8508 $
// SVN $Date: 2009-06-15 16:49:49 -0700 (Mon, 15 Jun 2009) $
`timescale 1ns/100ps
module
abfn_uart_1_sb_CoreUARTapb_0_0_fifo_256x8
(
CUARTI11
,
CUARTl11
,
CUARTOOOI
,
CUARTIOOI
,
WRB
,
RDB
,
RESET
,
FULL
,
EMPTY
)
;
output
[
7
:
0
]
CUARTI11
;
input
CUARTl11
;
input
CUARTOOOI
;
input
[
7
:
0
]
CUARTIOOI
;
input
WRB
;
input
RDB
;
input
RESET
;
output
FULL
;
output
EMPTY
;
parameter
[
6
:
0
]
CUARTIOlI
=
64
;
wire
[
7
:
0
]
CUARTI11
;
wire
AEMPTY
,
AFULL
,
FULL
,
EMPTY
;
abfn_uart_1_sb_CoreUARTapb_0_0_fifo_ctrl_128
CUARTIlOl
(
.CUARTOOII
(
CUARTIOOI
)
,
.CUARTIOII
(
CUARTI11
)
,
.CUARTOIlI
(
WRB
)
,
.CUARTIIlI
(
RDB
)
,
.CUARTlIlI
(
CUARTOOOI
)
,
.CUARTOllI
(
FULL
)
,
.CUARTIllI
(
EMPTY
)
,
.CUARTlllI
(
GEQTH
)
,
.CUARTlI
(
RESET
)
,
.CUARTIOlI
(
CUARTIOlI
)
)
;
endmodule
module
abfn_uart_1_sb_CoreUARTapb_0_0_fifo_ctrl_128
(
CUARTlIlI
,
CUARTlI
,
CUARTOOII
,
CUARTIIlI
,
CUARTOIlI
,
CUARTIOlI
,
CUARTIOII
,
CUARTOllI
,
CUARTIllI
,
CUARTlllI
)
;
parameter
CUARTO0lI
=
128
;
parameter
CUARTI0lI
=
7
;
parameter
CUARTl0lI
=
8
;
input
CUARTlIlI
;
input
CUARTlI
;
input
[
CUARTl0lI
-
1
:
0
]
CUARTOOII
;
input
CUARTIIlI
;
input
CUARTOIlI
;
input
[
6
:
0
]
CUARTIOlI
;
output
[
CUARTl0lI
-
1
:
0
]
CUARTIOII
;
output
CUARTOllI
;
output
CUARTIllI
;
output
CUARTlllI
;
wire
CUARTlIlI
;
wire
CUARTlI
;
wire
[
CUARTl0lI
-
1
:
0
]
CUARTOOII
;
wire
CUARTIIlI
;
wire
CUARTOIlI
;
reg
[
CUARTl0lI
-
1
:
0
]
CUARTIOII
;
wire
CUARTOllI
;
wire
CUARTIllI
;
wire
CUARTlllI
;
wire
[
CUARTl0lI
-
1
:
0
]
CUARTO1lI
;
reg
CUARTI1lI
;
reg
[
CUARTI0lI
-
1
:
0
]
CUARTl1lI
;
reg
[
CUARTI0lI
-
1
:
0
]
CUARTOO0I
;
reg
[
CUARTI0lI
-
1
:
0
]
CUARTIO0I
;
assign
CUARTOllI
=
(
CUARTl1lI
==
CUARTO0lI
-
1
)
?
1
'b
1
:
1
'b
0
;
assign
CUARTIllI
=
(
CUARTl1lI
==
0
)
?
1
'b
1
:
1
'b
0
;
assign
CUARTlllI
=
(
CUARTl1lI
>=
CUARTIOlI
)
?
1
'b
1
:
1
'b
0
;
always
@
(
posedge
CUARTlIlI
or
negedge
CUARTlI
)
begin
if
(
~
CUARTlI
)
begin
CUARTOO0I
<=
{
CUARTI0lI
{
1
'b
0
}
}
;
CUARTIO0I
<=
{
CUARTI0lI
{
1
'b
0
}
}
;
CUARTl1lI
<=
{
CUARTI0lI
{
1
'b
0
}
}
;
end
else
begin
if
(
~
CUARTIIlI
)
begin
if
(
CUARTOIlI
)
begin
CUARTl1lI
<=
CUARTl1lI
-
1
;
end
if
(
CUARTOO0I
==
CUARTO0lI
-
1
)
CUARTOO0I
<=
{
CUARTI0lI
{
1
'b
0
}
}
;
else
CUARTOO0I
<=
CUARTOO0I
+
1
;
end
if
(
~
CUARTOIlI
)
begin
if
(
CUARTl1lI
>=
CUARTO0lI
)
begin
$display
(
"\nERROR at time %0t:"
,
$time
)
;
$display
(
"FIFO Overflow\n"
)
;
$stop
;
end
if
(
CUARTIIlI
)
begin
CUARTl1lI
<=
CUARTl1lI
+
1
;
end
if
(
CUARTIO0I
==
CUARTO0lI
-
1
)
CUARTIO0I
<=
{
CUARTI0lI
{
1
'b
0
}
}
;
else
CUARTIO0I
<=
CUARTIO0I
+
1
;
end
end
end
always
@
(
posedge
CUARTlIlI
or
negedge
CUARTlI
)
begin
if
(
~
CUARTlI
)
begin
CUARTI1lI
<=
1
'b
0
;
CUARTIOII
<=
1
'b
0
;
end
else
begin
CUARTI1lI
<=
CUARTIIlI
;
if
(
CUARTI1lI
==
1
'b
0
)
begin
CUARTIOII
<=
CUARTO1lI
;
end
else
begin
CUARTIOII
<=
CUARTIOII
;
end
end
end
abfn_uart_1_sb_CoreUARTapb_0_0_ram128x8_pa4
CUARTllOl
(
.CUARTlO1I
(
CUARTOOII
)
,
.CUARTOI1I
(
CUARTO1lI
)
,
.CUARTII1I
(
CUARTIO0I
)
,
.CUARTlI1I
(
CUARTOO0I
)
,
.CUARTOl1I
(
CUARTOIlI
)
,
.CUARTll1I
(
CUARTlIlI
)
,
.CUARTO01I
(
CUARTlIlI
)
,
.CUARTlI
(
CUARTlI
)
)
;
endmodule
module
abfn_uart_1_sb_CoreUARTapb_0_0_ram128x8_pa4
(
CUARTlO1I
,
CUARTOI1I
,
CUARTII1I
,
CUARTlI1I
,
CUARTOl1I
,
CUARTll1I
,
CUARTO01I
,
CUARTlI
)
;
input
[
7
:
0
]
CUARTlO1I
;
input
[
6
:
0
]
CUARTII1I
,
CUARTlI1I
;
input
CUARTOl1I
,
CUARTll1I
,
CUARTO01I
,
CUARTlI
;
output
[
7
:
0
]
CUARTOI1I
;
wire
[
17
:
0
]
CUARTO0Ol
;
wire
CUARTl01I
,
VCC
,
GND
;
VCC
CUARTO11I
(
.Y
(
VCC
)
)
;
GND
CUARTI11I
(
.Y
(
GND
)
)
;
INV
CUARTl11I
(
.A
(
CUARTOl1I
)
,
.Y
(
CUARTl01I
)
)
;
assign
CUARTOI1I
=
CUARTO0Ol
[
7
:
0
]
;
RAM64x18
CUARTI0Ol
(
.A_DOUT
(
CUARTO0Ol
)
,
.B_DOUT
(
)
,
.BUSY
(
)
,
.A_ADDR_CLK
(
CUARTO01I
)
,
.A_DOUT_CLK
(
VCC
)
,
.A_ADDR_SRST_N
(
VCC
)
,
.A_DOUT_SRST_N
(
VCC
)
,
.A_ADDR_ARST_N
(
CUARTlI
)
,
.A_DOUT_ARST_N
(
VCC
)
,
.A_ADDR_EN
(
VCC
)
,
.A_DOUT_EN
(
VCC
)
,
.A_BLK
(
{
2
'b
11
}
)
,
.A_ADDR
(
{
CUARTlI1I
[
6
:
0
]
,
3
'b
0
}
)
,
.B_ADDR_CLK
(
VCC
)
,
.B_DOUT_CLK
(
VCC
)
,
.B_ADDR_SRST_N
(
VCC
)
,
.B_DOUT_SRST_N
(
VCC
)
,
.B_ADDR_ARST_N
(
VCC
)
,
.B_DOUT_ARST_N
(
VCC
)
,
.B_ADDR_EN
(
VCC
)
,
.B_DOUT_EN
(
VCC
)
,
.B_BLK
(
{
2
'b
0
}
)
,
.B_ADDR
(
{
10
'b
0
}
)
,
.C_CLK
(
CUARTll1I
)
,
.C_ADDR
(
{
CUARTII1I
[
6
:
0
]
,
3
'b
0
}
)
,
.C_DIN
(
{
10
'b
0
,
CUARTlO1I
[
7
:
0
]
}
)
,
.C_WEN
(
CUARTl01I
)
,
.C_BLK
(
{
2
'b
11
}
)
,
.A_EN
(
VCC
)
,
.A_ADDR_LAT
(
GND
)
,
.A_DOUT_LAT
(
VCC
)
,
.B_EN
(
GND
)
,
.B_ADDR_LAT
(
GND
)
,
.B_DOUT_LAT
(
VCC
)
,
.C_EN
(
VCC
)
,
.A_WIDTH
(
{
3
'b
011
}
)
,
.B_WIDTH
(
{
3
'b
011
}
)
,
.C_WIDTH
(
{
3
'b
011
}
)
,
.SII_LOCK
(
GND
)
)
;
endmodule
