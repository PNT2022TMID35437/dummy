//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Mon Aug 26 11:18:10 2024
// Version: 2024.1 2024.1.0.3
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// IIC
module IIC(
    // Inouts
    I2C_1_SCL,
    I2C_1_SDA
);

//--------------------------------------------------------------------
// Inout
//--------------------------------------------------------------------
inout  I2C_1_SCL;
inout  I2C_1_SDA;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   I2C_1_SCL;
wire   I2C_1_SDA;
wire   OSC_C0_0_RCOSC_25_50MHZ_O2F;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------IIC_MSS
IIC_MSS IIC_MSS_0(
        // Inputs
        .MCCC_CLK_BASE ( OSC_C0_0_RCOSC_25_50MHZ_O2F ),
        // Inouts
        .I2C_1_SDA     ( I2C_1_SDA ),
        .I2C_1_SCL     ( I2C_1_SCL ) 
        );

//--------OSC_C0
OSC_C0 OSC_C0_0(
        // Outputs
        .RCOSC_25_50MHZ_O2F ( OSC_C0_0_RCOSC_25_50MHZ_O2F ) 
        );


endmodule
